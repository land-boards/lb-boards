//���о΢����
//�绰 15815519071 QQ 906606596
//email : 906606596@qq.com 
//Email 906606596@qq.com
//ѧϰң�ؽ���������ԭ��
//�Ѱ��µļ�ͨ�������
//������ܵĵ�һλ��ʾ������ֵ�ķ���
//������ܵĵڶ�λ��ʾ������ֵ������
//�������Է�����λ����ܵ���ʾ�ǻ����ġ�
// learning remote control receiver decoding principle
//After pressing the key
//The first display keys complement digital tube
//Digital display of the second key key data
//You can find the results / two digital tube display is complementary.

module IR(clk,rst_n,IR,U2_138_select,U3_138_select,U2_138_A ,led_db);

  input   clk;  //ʱ������50M
  input   rst_n;
  input   IR;    //IR ����
  output [2:0] U2_138_A ;  //����138�ĵ�ַ������ܵ�λѡ�� 138 / control address, select the digital tube
  output [7:0] led_db;     //����ܵ����ݶ˿ڣ�/ / data port digital tube,
  output  U2_138_select;   //�����138ʹ�� Digital tube 138 enable
  output  U3_138_select;   //����138ʹ��  dot array 138 enable
 
  assign  U2_138_select = 1 ;  //ʹ�������138��Enable 138 digital tube, to make it work
  assign  U3_138_select = 0 ;  //�����õ���138������Will not let the dot array 138 work,
  reg [2:0] U2_138_A;
  reg [7:0] led_db;
 
  reg [7:0] led1,led2,led3,led4;
  reg [15:0] irda_data;    // save irda data,than send to 7 segment led
  reg [31:0] get_data;     // use for saving 32 bytes irda data
  reg [5:0]  data_cnt;     // 32 bytes irda data counter
  reg [2:0]  cs,ns;
  reg error_flag;          // 32 bytes data�ڼ䣬���ݴ����־

  //----------------------------------------------------------------------------
  reg irda_reg0;       //Ϊ�˱�������̬,������������Ĵ�������һ����ʹ�á�
  reg irda_reg1;       //����ſ���ʹ�ã����³����д���irda��״̬
  reg irda_reg2;       //Ϊ��ȷ��irda�ı��أ��ٴ�һ�μĴ��������³����д���irda��ǰһ״̬
  wire irda_neg_pulse; //ȷ��irda���½���
  wire irda_pos_pulse; //ȷ��irda��������
  wire irda_chang;     //ȷ�irda��������
  
  reg[15:0] cnt_scan;//ɨ��Ƶ�ʼ�����
   
  always @ (posedge clk) //�ڴ˲��ø���Ĵ���
    if(!rst_n)
      begin
        irda_reg0 <= 1'b0;
        irda_reg1 <= 1'b0;
        irda_reg2 <= 1'b0;
      end
    else
      begin
        irda_reg0 <= IR;
        irda_reg1 <= irda_reg0;
        irda_reg2 <= irda_reg1;
      end
     
  assign irda_chang = irda_neg_pulse | irda_pos_pulse;  //IR�����źŵĸı䣬���������½�
  assign irda_neg_pulse = irda_reg2 & (~irda_reg1);  //IR�����ź�irda�½���
  assign irda_pos_pulse = (~irda_reg2) & irda_reg1;      //IR�����ź�irda������

  //----------------------------------------------------------------------------
  //��Ʒ�Ƶ�ͼ������֣���PT2222�Ĺ淶�����Ƿ�����С�ĵ�ƽ���ʱ���?.56ms����
  //�����ڽ��в���ʱ��һ�㶼����ĵ�ƽ���?6�Ρ�Ҳ����˵Ҫ��0.56ms���ٲ���16
  //�Ρ�
  //              0.56ms/16=35us
  //?a href="javascript:;" onClick="javascript:tagshow(event, '%BF%AA%B7%A2');" 

//target="_self">���������Դ�����Ƶ?0MHz����ʱ������Ϊ20ns������������Ҫ�ķ�Ƶ����Ϊ��
  //              35000/20=1750
  //���������������������counter��һ��counter���ڼ�1750��ʱ����Ƶ��
  //һ��counter���ڼ����Ƶ֮��ͬһ�ֵ�ƽ��scan���ĵ���������������������ж�
  //��leader��9ms ����4.5ms���������ݵ� 0 ���� 1��
  //----------------------------------------------------------------------------
  reg [10:0] counter;  //��Ƶ1750��
  reg [8:0]  counter2; //������Ƶ��ĵ���
  wire check_9ms;  // check leader 9ms time
  wire check_4ms;  // check leader 4.5ms time
  wire low;        // check  data="0" time
  wire high;       // check  data="1" time
 
  //----------------------------------------------------------------------------
  //��Ƶ1750����
  always @ (posedge clk)
    if (!rst_n)
      counter <= 11'd0;
    else if (irda_chang)  //irda��ƽ�����ˣ������¿�ʼ����
      counter <= 11'd0;
    else if (counter == 11'd1750)
      counter <= 11'd0;
    else
      counter <= counter + 1'b1;
  
  //---------------------------------------------------------------------------- 
  always @ (posedge clk)
    if (!rst_n)
      counter2 <= 9'd0;
    else if (irda_chang)  //irda��ƽ�����ˣ������¿�ʼ�Ƶ�
      counter2 <= 9'd0;
    else if (counter == 11'd1750)
      counter2 <= counter2 +1'b1;
  

  assign check_9ms = ((217 < counter2) & (counter2 < 297)); 
  //257  Ϊ�������ȶ��ԣ�ȡһ����Χ
  assign check_4ms = ((88 < counter2) & (counter2 < 168));  //128
  assign low  = ((6 < counter2) & (counter2 < 26));         // 16
  assign high = ((38 < counter2) & (counter2 < 58));        // 48

  //----------------------------------------------------------------------------
  // generate statemachine  ״̬��
    parameter IDLE       = 3'b000, //��ʼ״̬
              LEADER_9   = 3'b001, //9ms
              LEADER_4   = 3'b010, //4ms
              DATA_STATE = 3'b100; //��������
 
  always @ (posedge clk)
    if (!rst_n)
      cs <= IDLE;
    else
      cs <= ns; //״̬λ
     
  always @ ( * )
    case (cs)
      IDLE:
        if (~irda_reg1)
          ns = LEADER_9;
        else
          ns = IDLE;
   
      LEADER_9:
        if (irda_pos_pulse)   //leader 9ms check
          begin
            if (check_9ms)
              ns = LEADER_4;
            else
              ns = IDLE;
          end
        else  //�걸��if---else--- ;��ֹ����latch
          ns =LEADER_9;
   
      LEADER_4:
        if (irda_neg_pulse)  // leader 4.5ms check
          begin
            if (check_4ms)
              ns = DATA_STATE;
            else
              ns = IDLE;
          end
        else
          ns = LEADER_4;
   
      DATA_STATE:
        if ((data_cnt == 6'd32) & irda_reg2 & irda_reg1)
          ns = IDLE;
        else if (error_flag)
          ns = IDLE;
        else
          ns = DATA_STATE;
      default:
        ns = IDLE;
    endcase

  //״̬���е����,��ʱ���·������
  always @ (posedge clk)
    if (!rst_n)
      begin
        data_cnt <= 6'd0;
        get_data <= 32'd0;
        error_flag <= 1'b0;
      end
  
    else if (cs == IDLE)
      begin
        data_cnt <= 6'd0;
        get_data <= 32'd0; 
        error_flag <= 1'b0;
      end
  
    else if (cs == DATA_STATE)
      begin
        if (irda_pos_pulse)  // low 0.56ms check
          begin
            if (!low)  //error
              error_flag <= 1'b1;
          end
        else if (irda_neg_pulse)  //check 0.56ms/1.68ms data 0/1
          begin
            if (low)
              get_data[0] <= 1'b0;
            else if (high)
              get_data[0] <= 1'b1;
            else
              error_flag <= 1'b1;
             
            get_data[31:1] <= get_data[30:0];
            data_cnt <= data_cnt + 1'b1;
          end
      end

  always @ (posedge clk)
    if (!rst_n)
      irda_data <= 16'd0;
    else if ((data_cnt ==6'd32) & irda_reg1)
  begin
   led1 <= get_data[7:0];  //���ݷ���
   led2 <= get_data[15:8]; //������
   led3 <= get_data[23:16];//�û���
   led4 <= get_data[31:24];
  end
 
 //�����ɨ���õ��ļ�����
always@(posedge clk or negedge  rst_n)
begin
	if(!rst_n) begin
		cnt_scan<=0;
		
	 end
	else begin
		cnt_scan<=cnt_scan+1;
		end
end
//��λ����ܵõ�������ʾ��ʱ��
always @(cnt_scan)
begin
   case(cnt_scan[15:14])
       2'b00 :
          U2_138_A = 3'b000;  
       2'b01 :
          U2_138_A = 3'b001;
   //    2'b10 :
    //      led_cs = 4'b1011;
    //   2'b11 :
   //       led_cs = 4'b0111;
       default :
          U2_138_A = 3'b000;
    endcase
end

//�û���Ҫע�⣬������ʾ����ң�ذ�ÿһ�������ı���ֵ��
//������˵���Ұ���һ��1�� ������ʾ1������ʾ��1�ⰴ�����롣
//����ÿ������һ�����֤һ���ģ�
always@(U2_138_A) 
begin
	case(U2_138_A)
		3'b000:
			led_db<= led1; //������ܵĵ�һλ��ʾ������ֵ�ķ���
		3'b001:
			led_db<= led2; //������ܵĵڶ�λ��ʾ������ֵ������
	//	4'b1011:
	//		led_db<= led3;
	//	4'b0111:
	//		led_db<= led4;
	  

	 endcase
end

endmodule 


